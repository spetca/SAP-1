module output_reg(
    input [7:0] dbus, 
    input n_lo, 
    input clk, 
    output [7:0] bdisp
);

endmodule